module Rcon(i,rcon);
input [3:0]i;
output [31:0] rcon;

assign rcon=(i== 4'd0)?32'h01_00_00_00:
      (i==   4'd1)? 32'h02_00_00_00:
         (i==4'd2)? 32'h04_00_00_00:
       (i==  4'd3)?32'h08_00_00_00:
        (i== 4'd4)?32'h10_00_00_00:
        (i== 4'd5)?32'h20_00_00_00:
        (i== 4'd6)?32'h40_00_00_00:
         (i==4'd7) ?32'h80_00_00_00:
         (i==4'd8)?32'h1b_00_00_00:
       (i==  4'd9) ?32'h36_00_00_00:
			(i==4'd10) ?32'h6C_00_00_00:
			(i==4'd11) ?32'hD8_00_00_00:
			(i==4'd12) ?32'h23_00_00_00:
			(i==4'd13)	?32'h46_00_00_00:0;
		
			
        


endmodule